module phase_to_angle_converter(
  input       reset,
  input [N:0] phase_in,     // Phase input
  input [N:0] amplitude_in, // Amplitude input
  
  output reg [2*N:0] out      // Angle output
);

parameter N = 8;

reg [N:0] LUT [0:511];

initial
begin
    LUT[0] = 256;
	LUT[1] = 259;
	LUT[2] = 262;
	LUT[3] = 265;
	LUT[4] = 269;
	LUT[5] = 272;
	LUT[6] = 275;
	LUT[7] = 278;
	LUT[8] = 281;
	LUT[9] = 284;
	LUT[10] = 287;
	LUT[11] = 290;
	LUT[12] = 294;
	LUT[13] = 297;
	LUT[14] = 300;
	LUT[15] = 303;
	LUT[16] = 306;
	LUT[17] = 309;
	LUT[18] = 312;
	LUT[19] = 315;
	LUT[20] = 318;
	LUT[21] = 321;
	LUT[22] = 324;
	LUT[23] = 327;
	LUT[24] = 330;
	LUT[25] = 333;
	LUT[26] = 336;
	LUT[27] = 339;
	LUT[28] = 342;
	LUT[29] = 345;
	LUT[30] = 348;
	LUT[31] = 351;
	LUT[32] = 354;
	LUT[33] = 357;
	LUT[34] = 360;
	LUT[35] = 363;
	LUT[36] = 365;
	LUT[37] = 368;
	LUT[38] = 371;
	LUT[39] = 374;
	LUT[40] = 377;
	LUT[41] = 379;
	LUT[42] = 382;
	LUT[43] = 385;
	LUT[44] = 388;
	LUT[45] = 390;
	LUT[46] = 393;
	LUT[47] = 396;
	LUT[48] = 398;
	LUT[49] = 401;
	LUT[50] = 403;
	LUT[51] = 406;
	LUT[52] = 408;
	LUT[53] = 411;
	LUT[54] = 413;
	LUT[55] = 416;
	LUT[56] = 418;
	LUT[57] = 421;
	LUT[58] = 423;
	LUT[59] = 426;
	LUT[60] = 428;
	LUT[61] = 430;
	LUT[62] = 433;
	LUT[63] = 435;
	LUT[64] = 437;
	LUT[65] = 439;
	LUT[66] = 441;
	LUT[67] = 444;
	LUT[68] = 446;
	LUT[69] = 448;
	LUT[70] = 450;
	LUT[71] = 452;
	LUT[72] = 454;
	LUT[73] = 456;
	LUT[74] = 458;
	LUT[75] = 460;
	LUT[76] = 462;
	LUT[77] = 463;
	LUT[78] = 465;
	LUT[79] = 467;
	LUT[80] = 469;
	LUT[81] = 471;
	LUT[82] = 472;
	LUT[83] = 474;
	LUT[84] = 476;
	LUT[85] = 477;
	LUT[86] = 479;
	LUT[87] = 480;
	LUT[88] = 482;
	LUT[89] = 483;
	LUT[90] = 485;
	LUT[91] = 486;
	LUT[92] = 487;
	LUT[93] = 489;
	LUT[94] = 490;
	LUT[95] = 491;
	LUT[96] = 493;
	LUT[97] = 494;
	LUT[98] = 495;
	LUT[99] = 496;
	LUT[100] = 497;
	LUT[101] = 498;
	LUT[102] = 499;
	LUT[103] = 500;
	LUT[104] = 501;
	LUT[105] = 502;
	LUT[106] = 503;
	LUT[107] = 504;
	LUT[108] = 504;
	LUT[109] = 505;
	LUT[110] = 506;
	LUT[111] = 506;
	LUT[112] = 507;
	LUT[113] = 508;
	LUT[114] = 508;
	LUT[115] = 509;
	LUT[116] = 509;
	LUT[117] = 510;
	LUT[118] = 510;
	LUT[119] = 510;
	LUT[120] = 511;
	LUT[121] = 511;
	LUT[122] = 511;
	LUT[123] = 511;
	LUT[124] = 511;
	LUT[125] = 511;
	LUT[126] = 511;
	LUT[127] = 511;
	LUT[128] = 511;
	LUT[129] = 511;
	LUT[130] = 511;
	LUT[131] = 511;
	LUT[132] = 511;
	LUT[133] = 511;
	LUT[134] = 511;
	LUT[135] = 511;
	LUT[136] = 511;
	LUT[137] = 510;
	LUT[138] = 510;
	LUT[139] = 510;
	LUT[140] = 509;
	LUT[141] = 509;
	LUT[142] = 508;
	LUT[143] = 508;
	LUT[144] = 507;
	LUT[145] = 506;
	LUT[146] = 506;
	LUT[147] = 505;
	LUT[148] = 504;
	LUT[149] = 504;
	LUT[150] = 503;
	LUT[151] = 502;
	LUT[152] = 501;
	LUT[153] = 500;
	LUT[154] = 499;
	LUT[155] = 498;
	LUT[156] = 497;
	LUT[157] = 496;
	LUT[158] = 495;
	LUT[159] = 494;
	LUT[160] = 493;
	LUT[161] = 491;
	LUT[162] = 490;
	LUT[163] = 489;
	LUT[164] = 487;
	LUT[165] = 486;
	LUT[166] = 485;
	LUT[167] = 483;
	LUT[168] = 482;
	LUT[169] = 480;
	LUT[170] = 479;
	LUT[171] = 477;
	LUT[172] = 476;
	LUT[173] = 474;
	LUT[174] = 472;
	LUT[175] = 471;
	LUT[176] = 469;
	LUT[177] = 467;
	LUT[178] = 465;
	LUT[179] = 463;
	LUT[180] = 462;
	LUT[181] = 460;
	LUT[182] = 458;
	LUT[183] = 456;
	LUT[184] = 454;
	LUT[185] = 452;
	LUT[186] = 450;
	LUT[187] = 448;
	LUT[188] = 446;
	LUT[189] = 444;
	LUT[190] = 441;
	LUT[191] = 439;
	LUT[192] = 437;
	LUT[193] = 435;
	LUT[194] = 433;
	LUT[195] = 430;
	LUT[196] = 428;
	LUT[197] = 426;
	LUT[198] = 423;
	LUT[199] = 421;
	LUT[200] = 418;
	LUT[201] = 416;
	LUT[202] = 413;
	LUT[203] = 411;
	LUT[204] = 408;
	LUT[205] = 406;
	LUT[206] = 403;
	LUT[207] = 401;
	LUT[208] = 398;
	LUT[209] = 396;
	LUT[210] = 393;
	LUT[211] = 390;
	LUT[212] = 388;
	LUT[213] = 385;
	LUT[214] = 382;
	LUT[215] = 379;
	LUT[216] = 377;
	LUT[217] = 374;
	LUT[218] = 371;
	LUT[219] = 368;
	LUT[220] = 365;
	LUT[221] = 363;
	LUT[222] = 360;
	LUT[223] = 357;
	LUT[224] = 354;
	LUT[225] = 351;
	LUT[226] = 348;
	LUT[227] = 345;
	LUT[228] = 342;
	LUT[229] = 339;
	LUT[230] = 336;
	LUT[231] = 333;
	LUT[232] = 330;
	LUT[233] = 327;
	LUT[234] = 324;
	LUT[235] = 321;
	LUT[236] = 318;
	LUT[237] = 315;
	LUT[238] = 312;
	LUT[239] = 309;
	LUT[240] = 306;
	LUT[241] = 303;
	LUT[242] = 300;
	LUT[243] = 297;
	LUT[244] = 294;
	LUT[245] = 290;
	LUT[246] = 287;
	LUT[247] = 284;
	LUT[248] = 281;
	LUT[249] = 278;
	LUT[250] = 275;
	LUT[251] = 272;
	LUT[252] = 269;
	LUT[253] = 265;
	LUT[254] = 262;
	LUT[255] = 259;
	LUT[256] = 256;
	LUT[257] = 253;
	LUT[258] = 250;
	LUT[259] = 247;
	LUT[260] = 243;
	LUT[261] = 240;
	LUT[262] = 237;
	LUT[263] = 234;
	LUT[264] = 231;
	LUT[265] = 228;
	LUT[266] = 225;
	LUT[267] = 222;
	LUT[268] = 218;
	LUT[269] = 215;
	LUT[270] = 212;
	LUT[271] = 209;
	LUT[272] = 206;
	LUT[273] = 203;
	LUT[274] = 200;
	LUT[275] = 197;
	LUT[276] = 194;
	LUT[277] = 191;
	LUT[278] = 188;
	LUT[279] = 185;
	LUT[280] = 182;
	LUT[281] = 179;
	LUT[282] = 176;
	LUT[283] = 173;
	LUT[284] = 170;
	LUT[285] = 167;
	LUT[286] = 164;
	LUT[287] = 161;
	LUT[288] = 158;
	LUT[289] = 155;
	LUT[290] = 152;
	LUT[291] = 149;
	LUT[292] = 147;
	LUT[293] = 144;
	LUT[294] = 141;
	LUT[295] = 138;
	LUT[296] = 135;
	LUT[297] = 133;
	LUT[298] = 130;
	LUT[299] = 127;
	LUT[300] = 124;
	LUT[301] = 122;
	LUT[302] = 119;
	LUT[303] = 116;
	LUT[304] = 114;
	LUT[305] = 111;
	LUT[306] = 109;
	LUT[307] = 106;
	LUT[308] = 104;
	LUT[309] = 101;
	LUT[310] = 99;
	LUT[311] = 96;
	LUT[312] = 94;
	LUT[313] = 91;
	LUT[314] = 89;
	LUT[315] = 86;
	LUT[316] = 84;
	LUT[317] = 82;
	LUT[318] = 79;
	LUT[319] = 77;
	LUT[320] = 75;
	LUT[321] = 73;
	LUT[322] = 71;
	LUT[323] = 68;
	LUT[324] = 66;
	LUT[325] = 64;
	LUT[326] = 62;
	LUT[327] = 60;
	LUT[328] = 58;
	LUT[329] = 56;
	LUT[330] = 54;
	LUT[331] = 52;
	LUT[332] = 50;
	LUT[333] = 49;
	LUT[334] = 47;
	LUT[335] = 45;
	LUT[336] = 43;
	LUT[337] = 41;
	LUT[338] = 40;
	LUT[339] = 38;
	LUT[340] = 36;
	LUT[341] = 35;
	LUT[342] = 33;
	LUT[343] = 32;
	LUT[344] = 30;
	LUT[345] = 29;
	LUT[346] = 27;
	LUT[347] = 26;
	LUT[348] = 25;
	LUT[349] = 23;
	LUT[350] = 22;
	LUT[351] = 21;
	LUT[352] = 19;
	LUT[353] = 18;
	LUT[354] = 17;
	LUT[355] = 16;
	LUT[356] = 15;
	LUT[357] = 14;
	LUT[358] = 13;
	LUT[359] = 12;
	LUT[360] = 11;
	LUT[361] = 10;
	LUT[362] = 9;
	LUT[363] = 8;
	LUT[364] = 8;
	LUT[365] = 7;
	LUT[366] = 6;
	LUT[367] = 6;
	LUT[368] = 5;
	LUT[369] = 4;
	LUT[370] = 4;
	LUT[371] = 3;
	LUT[372] = 3;
	LUT[373] = 2;
	LUT[374] = 2;
	LUT[375] = 2;
	LUT[376] = 1;
	LUT[377] = 1;
	LUT[378] = 1;
	LUT[379] = 0;
	LUT[380] = 0;
	LUT[381] = 0;
	LUT[382] = 0;
	LUT[383] = 0;
	LUT[384] = 0;
	LUT[385] = 0;
	LUT[386] = 0;
	LUT[387] = 0;
	LUT[388] = 0;
	LUT[389] = 0;
	LUT[390] = 1;
	LUT[391] = 1;
	LUT[392] = 1;
	LUT[393] = 2;
	LUT[394] = 2;
	LUT[395] = 2;
	LUT[396] = 3;
	LUT[397] = 3;
	LUT[398] = 4;
	LUT[399] = 4;
	LUT[400] = 5;
	LUT[401] = 6;
	LUT[402] = 6;
	LUT[403] = 7;
	LUT[404] = 8;
	LUT[405] = 8;
	LUT[406] = 9;
	LUT[407] = 10;
	LUT[408] = 11;
	LUT[409] = 12;
	LUT[410] = 13;
	LUT[411] = 14;
	LUT[412] = 15;
	LUT[413] = 16;
	LUT[414] = 17;
	LUT[415] = 18;
	LUT[416] = 19;
	LUT[417] = 21;
	LUT[418] = 22;
	LUT[419] = 23;
	LUT[420] = 25;
	LUT[421] = 26;
	LUT[422] = 27;
	LUT[423] = 29;
	LUT[424] = 30;
	LUT[425] = 32;
	LUT[426] = 33;
	LUT[427] = 35;
	LUT[428] = 36;
	LUT[429] = 38;
	LUT[430] = 40;
	LUT[431] = 41;
	LUT[432] = 43;
	LUT[433] = 45;
	LUT[434] = 47;
	LUT[435] = 49;
	LUT[436] = 50;
	LUT[437] = 52;
	LUT[438] = 54;
	LUT[439] = 56;
	LUT[440] = 58;
	LUT[441] = 60;
	LUT[442] = 62;
	LUT[443] = 64;
	LUT[444] = 66;
	LUT[445] = 68;
	LUT[446] = 71;
	LUT[447] = 73;
	LUT[448] = 75;
	LUT[449] = 77;
	LUT[450] = 79;
	LUT[451] = 82;
	LUT[452] = 84;
	LUT[453] = 86;
	LUT[454] = 89;
	LUT[455] = 91;
	LUT[456] = 94;
	LUT[457] = 96;
	LUT[458] = 99;
	LUT[459] = 101;
	LUT[460] = 104;
	LUT[461] = 106;
	LUT[462] = 109;
	LUT[463] = 111;
	LUT[464] = 114;
	LUT[465] = 116;
	LUT[466] = 119;
	LUT[467] = 122;
	LUT[468] = 124;
	LUT[469] = 127;
	LUT[470] = 130;
	LUT[471] = 133;
	LUT[472] = 135;
	LUT[473] = 138;
	LUT[474] = 141;
	LUT[475] = 144;
	LUT[476] = 147;
	LUT[477] = 149;
	LUT[478] = 152;
	LUT[479] = 155;
	LUT[480] = 158;
	LUT[481] = 161;
	LUT[482] = 164;
	LUT[483] = 167;
	LUT[484] = 170;
	LUT[485] = 173;
	LUT[486] = 176;
	LUT[487] = 179;
	LUT[488] = 182;
	LUT[489] = 185;
	LUT[490] = 188;
	LUT[491] = 191;
	LUT[492] = 194;
	LUT[493] = 197;
	LUT[494] = 200;
	LUT[495] = 203;
	LUT[496] = 206;
	LUT[497] = 209;
	LUT[498] = 212;
	LUT[499] = 215;
	LUT[500] = 218;
	LUT[501] = 222;
	LUT[502] = 225;
	LUT[503] = 228;
	LUT[504] = 231;
	LUT[505] = 234;
	LUT[506] = 237;
	LUT[507] = 240;
	LUT[508] = 243;
	LUT[509] = 247;
	LUT[510] = 250;
	LUT[511] = 253;
end

always @(posedge reset)
begin
out <= 0;
end

always @(*) 
begin
  out = LUT[phase_in] * amplitude_in;
  //$readmemh("lut.txt", LUT);
end

endmodule


/*
	Our tiny RISC-V CPU
*/
module cpurv(
	input clock,
	input reset,
	
	output [31:0] progaddress,
	input  [31:0] instruction,
	
	output [31:0] dataoutport,
	input  [31:0] datainport
	);

// Local wires:

wire [ 1:0] pcfunc;  // function to define the next value of PC (2 bits)
			            // 00: PC<=PC+4;  
					      // 01: PC<=PC+immediate;
					     	// 10: PC<=PC+rs1+immediate
					     	// 11: PC<=PC+immediate<<12

wire [21:0] pcoffset;   // signed offset to add to PC (22 bits)

wire [31:0] pcaddress;  // the current value of program counter (32 bits)

wire [31:0] regdatain;    // input data to write in the register specified by writeselect[4:0]

wire [ 4:0] readselect1, readselect2, writeselect; // read and write register selectors

wire        writeenable;  // enable writting to a register

wire [31:0] regdataout1, regdataout2;  // The output data from the register file, goes to the ALU

wire [31:0] dataimmed;    // Immediate data deoced from the intruction to the ALU

wire        selopr2;      // Select the 2nd operand to the ALU: 0=rdatain2, 1=dataimmed

wire [ 3:0] aluoper;	  // ALU operation, must be coherent between the decoder and the ALU impltation

wire [31:0] aluresult;    // The result generated by the ALU, 32 bits

wire        aluzeroflag;  // Zero flag: is 1 if current result is zero.

//--------------------------------------------------------------------------------- 	
// The program counter (PC) logic:
programcounter programcounter_1
          (
		    .clock( clock ),
			.reset( reset ),	
			.func(  pcfunc ),       // function to define the next value of PC (2 bits)
			                        // 00: PC<=PC+4;  
								    // 01: PC<=PC+immediate;
								    // 10: PC<=PC+rs1+immediate
								    // 11: PC<=PC+immediate<<12
								  
			.offset( pcoffset ),    // signed offset to add to PC (22 bits) -- immediate
						
			.rs1( readselect1 ),    // read select 1, 5 bits (0 .. 31)
			
			.pcout( pcaddress )  // the current value of PC (32 bits)
		  );

//---------------------------------------------------------------------------------                   	
// The register file logic: 32 registers, 32-bit names x0 to x31
// register x0 is readonly and always returns zero.
regfile regfile_1
           (
		     .clock( clock ),
			 .reset( reset ),
			 .datain( regdatain ),		// datain to write into a register, 32 bits
			 .rs1( readselect1 ),		// read select 1, 5 bits (0 .. 31)
			 .rs2( readselect2 ),		// read select 2, 5 bits (0 .. 31)
			 .we( writeenable ),        // write enable, set to 1 to write regdatain into register writeselect
			 .rd( writeselect ),        // index of register to write, 5 bits, (0..31)
			 .dataout1( regdataout1 ),  // data out 1, contents of register selected by rs1
			 .dataout2( regdataout2 )   // data out 2, contents of register selected by rs2
		   );

//---------------------------------------------------------------------------------		   
// The ALU: implements up to 16 operations specf'd by aluoper
// two 32-bit inputs, one 32-bit output, one 1-bit output (zero flag)
alu  alu_1
			(
			  .clock( clock ),
			  .reset( reset ),
			  .rdatain1( regdataout1 ),	// operand 1 (rs1), 32 bits
			  .rdatain2( regdataout2 ),	// operand 2 (rs2), 32 bits
			  .dataimmed( dataimmed ),  // immediate data in, 32 bits
			  .selopr2( selopr2 ),      // Select the 2nd operand to the ALU: 0=rdatain2, 1=dataimmed
			  .aluoper( aluoper ),      // ALU operation, 4 bits
			  .aluresult( aluresult ),	// result of the ALU operation, 32 bits
			  .zero( aluzeroflag )
			);

//---------------------------------------------------------------------------------
// Instruction decoder: receives the 32-bit instruction and generates
// the various control signals:
decodeinstruction decodeinstruction_1
			(
			  .instruction( instruction ),  // The instruction read from the program memory
			  
			  // control of program counter:
			  .pcfunc( pcfunc ),			// 2-bit function for PC update (see above)
			  .pcoffset( pcoffset ),		// the immediate data extracted from the instruction 
			                                // to add to the PC, in the case of branch instructions
			                                
			  
			  // control of the register file:
			  .readselect1( readselect1 ),  // read select for operand rs1
			  .readselect2( readselect2 ),  // read select for operand rs2
			  .writeenable( writeenable ),  // write enable 
			  .writeselect( writeselect ),  // Index of register to write
			  
			  // control of the ALU:
			  .aluoper( aluoper ),			// ALU operation, 4 bits, up to 16 operations
			  .selopr2( selopr2 ),			// Select the 2nd operand to the ALU: 0=rdatain2, 1=dataimmed
			  
			  // immediate data:
			  .immediate( dataimmed )		// immediate data for the 2nd operand of the ALU, 32 bits.
			                                // Note that some immediates extracted from the instructions
											// are shorter than 32 bits but must be extended to 32 bits
											// to enter the ALU 2nd operand
			);

// Local connections:
// This version does not support data memory instructions
// ALU result is connected directly to the datain port of the register file:
assign regdatain = aluresult;
	
endmodule	
	
	
